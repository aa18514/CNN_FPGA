XlxV61EB    2999     8b0a	��UV�.��=�@���}t[���A�u{�wZ�}�?
g]H2:�n�.�d��:S� \`?D��>s<X�@sRZ�%��P$R�	a�'|��Ď��NWuӀ���$�Of9ڲ�Jm쇪����ņ|�l50ٸF�;�ͦY4nm8Q��������s��/�GչQEN7T��]��8���Z�ȹi%ky5�]>�-��w0H:��uo����=6�������Z�NX��?�d'�^`�.�1\��#�~T�d|��.��-N ��Ѵh�m������)5�<B}R�;`�9��(��3� �b�?�{p� <
�F�-w�]��:ƴ �n�~��ĉ�Ly��g-l`[��n4�f(b�-ܽ�����@{�E�[1���98i�Mha ����] �g�	l{q����+FN����]g��`\a@έ� ��n�!>.�;��໓��D�'�a���Zu� %0�Q�Ef�|��d����S����':q�v߃V�g����!��&pR���E�'JsA30�Z�-wpwZ[.�z4ŵ�>�0�Ո���Z��@}*5C�%��Ȃkz	��v��=����՞_f�&`a�ߒ�j\���Z�>�����Y�G���\]Kr:�~O���X�c���7��~@ ��5�lX4��`���k�&�2������q:��]5{�:�tB�2I�⬑|�D��܏��ҙI�^7m�'t: �1���M�����]^�_�įs���i"��@�M'h�k橵�s�F˄�Ѿ�[	��߸���M`��_[������*����)Vs�|�Y�s��$��!�(����|�[�_�������+#K�`Ҧ?uc=�Ԗ9�o�֎��^�yݳ	�`!ƃ��m�A�&���#��&��ßi�MvJʃ	9�y}P*A��nx4U=`�?�F���Q�ᅯ��	���{p�OU�5�Y��U��h�qN��[;��ʖ-���c��<�
��$�
�m�P	
-��V <���ޔ��ގﮃ"O�&䶾"8L�(���-ptK�9%�����>��;����k�;!ot�O���zT�ϼ��y���u[e�Ӧ."Ӑ���,Ɗ� �Y����%�i�/� 'o쿮����.��(N$y?�h�P��U(O��4���|p*�a1���9/L�Y-�j6�6~Z$�/�j���)P�7%�l����W���0@Mߍтd��[y� �����T�Ȇ�k�ѣb<�{��s.#����NÇ����=���L�#�M#��»#�6͵A������E����N���ev��|�>4ː ����@�ϗ�Iҵ��)�0��:^�C~'нuc�U�j6������a+~!�.B�-Ry��2"zu�?O,�	�#�I�"��X݈�O"��iɷǦ��.��Z�H�~V�s�����}!�:���Co{��<�r��M=}�_u��=���Ұ��$G�V�-���g8���̪���M�S�Zz�yx��+���~�����O�捴�C=�M� ^(�{���{q���j��=�ҁ��m��7����t<N4t��1TK��3J>P����)�E�<����OE��e��
��L�g��.�����:��z��Lπ���!|�
˜�2"Y���A�5p�{j���#�'"�����ֆ鳪1P�0��p����a�EH�z�9�b������"�Nu����>B�����7s���7�d���x
]���S�io;��[q~���)�c⠽x�>~1,]2�W��d,hRׯ�N��C3�T-�c_�6�e$O�Хh:��
��9lW�j��dU��i�b���a|�9��'�WF��Q'���S'y|���uL�<���6h��G	a�T����|�����P~��c���E�|Z(y_r�>��5s�����Q����O.�&�l�E���D��J�Ѽۘ��S:�F�� �%���0��������ײ��)>"a�iDq3B���(���$��s�+%S)��Wٮ��+bًM�$����m��&4�Tt����N�zP�V{��D9�T��]���uR>i,�Cw���X���fG~"T�[�6�yj�CK'፛��ᢌ���"��)5����>|]��Y�0�sj�V`?��g��j��