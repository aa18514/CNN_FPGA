XlxV61EB    1cbe     7f0��=�^iq�ѯ���3��r���jH�.jj)�I=����ua55�!�1��)��3��O��)�Da��Y^$[�Mƣ���QO'1���<ɟ�w��3�5ۖ5 ��N�¦�e���k؂��ji̍��B�l��G����l$Y��9s��8�t�{x/2��~Ӑ~��?���Ll;]��-#���L4��C�i$� � ��yO��G!�[B���P��\n },c��}���Ɵ�[�Ta�ߤ�dA�	3��-��<d��rF��m	�\�':���2#6���V��"8_���N�/�%�t��~��[�㭚��Y��p+]|:Z�y�U�ſ8�M����I�=�T)������ۤ�^|Ƙ>��<*z�z=**7��)^d�̙z2��J��	��61��c0}Q��N�T����8��@�;�o�3��3M�ύ�p�a/6��^���+8a�I]�J�Q4����$'3��x�����x���@��5J>����.��*�"ZO���o���{t�8�GP�6�.�W��0� v��
&��� �-����92&24�N�X�}~���X���Т�!�X�k�&	eg��T�\M�pEĞ��� G`��l�|�6�P�Gƛٌ���V򝞅��N�,�w���O{�|=C{x7��qD�kJ�2�QA�}�9�$x��"J�B>���M��׬��Y�ւt�P1=����u�}��)ﲜ��b��L�ʊ@�`�i�.��B���4Tc	�CT��RԾ:)�s` �?�i!�Β��1�������B7��FmH-s�`��J׵�ȪN�ل�z)(^l��fD����(=+U�=rKK�=�8@~����3ET���*[���<5|&7N2j���S��"�g@���wS>�E��A���~���2��1T����e�a� ���l�M���>=r���/�bc���	�D<d�:��H��E$f]����:ڮ,��f�S�y(e��O{QՔ*��	�Ri�]�AZ�9J����G\��sˮ��~^
Hj(S�x����ѝc�P��u_�~O��У�{�֐��2S�����ps� /�dm#��5@z���4�HJ�cGnԢʝ§��2�_=��Hi%~�E�~��d�OX��� ��-�;�/R��݌�2���L�rǁP7,+Rc�9A���"�D��L�T�~a����u���,t!�9ʈ�I�̟f]����3�6�<B(>�=��+h�L+k��	iV�gr!8c� i ߘ����n?H��c|So~.�J��9z�p	�*��
X"٩#�dP�}�"Z����Y���r��������Y��Ѳ� X^:�� ��[^g��u�k1g-`MǡJ+����`�i=-�K�CP��kAye����?$N�wΫ�j�:I�*�a ���~�g�es���'*x�~*y$�G�(��>ͫˎ����`wbF�I�-��>ڢ�Q��\Q�����XA�Z��A�),����V�5k\Ä��Z!������_�!< �4q��`�z�5!ix�dr��	���):� |��.���[DV���B�d9]�h�>ȚbO9����{����H��\$j��� ;N7(
Z��)���ڸ��hݐЖW������ȡif�4�E��.܋���)��1;;Q���ޑ˱���a8ǭ�xW����AA�'�v�(��v�*���,��0$ý�B�Pc��XQ�L 1����~  �%x�8O�4���3�5�u�R5���M��u1ثa>�ϛUr4�űT���ѵ�.�FbO͎������>�Ԙ��KlSC،7���ri�n3"::��^ #"n'h�e�^��|�"�>+E�`j�#p������Z�@� �gkh�FV}ݫ��k�}|D6/�K�0�1�Q!�h��p�Rf�,�\5�;iB_�h'��h�)Re�'��I�1e.^l�Rk<�T�jNd�D��3*��a[D}ͮ]|�����Ÿ���R���U��Ѷ ���2����g