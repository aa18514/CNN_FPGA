XlxV61EB    5258    1260���̋L����o�rwx��m�vQd�j�H�$�w��=#3�6�r����l]?-���d'�"�l�N��l��=�塜���+m���O0=�Wh���XI�=D	�I�=���U��Rx���<ge��|�o�;�����������>y_��8�+�=� �}R6�K?�f'�6�sȃ�N����SY�:��H�m�2țb6�S#�]X��}��%W~��6��\�a)/n�>���v�oP\*;8��R6���!
5-;wƜ=L3i?Z'��F�2�>)�!�y���'+����ƈ��v�V�C~�ڙ��F��(V���w/$�S]���\���|�E[q�V�<wi@�`���)��j����pT�]�O�/"dP6��5.��)M����ʍf��Ù_��f(��|��"�7÷��JYF����B!	�+p��r�)�sORYk4����ؚ᫆/�Y��hI��~1���Ghjg�e��Z�O���Z��[4r/��ޘi̱Y-aZ�#��MM���`I�+"�&!�Kz�8���"-�Д�c�¢�=8��1��	|��O\��d��(��sw0`�l\Q+S�!Z�"�OST�ǣ�-~P��8��>�\���2�9]�
�0t�cw.�9��|
�L���"���ݜ��'z�8m���5r����WX@��i�	���R>����!��:C��Z��:��j��k��s�G�'eo��L�>��˖r�s.�2��V�ikv Pd:$�B�Ys�	��P���e�0ovNF��JXň�+���܁v��}�"�C"���|X��-i��Z���ur�Z ]�gəĚ�7e���9�VX�LI���t�(��!���~�3���K�U;�����$TR��;	���N�Ŭ��̀ 	�MVU7}&��(��� ֡�}�����9cӶe�.UX�yؖF� ��_�%n�L����?;YF��dUҦ����	ʭ0���o%-��&�'�b]4O�wi���8���t�c�Rb�a9�1[ %��b��^|���䞬��UFj��\B~��ӗ�	�� 7�IF�w�kyuHÛ�j�A�J`���6����Q���'�,� �S�V3\.����g�6���s/sCOG��zA��o1���A�������^��\��9,r!bA�iZ֘�Ƈ�Yu|9*���ѭ�n0�/�
���u�Rx����_�g�D�2�Q�,��N��;����#B�p&�~��2l5��n��c:ǟF�^��#�3A�]��"� �NC,w�����	g��BBO_,?O�����>5ʏ�=�Ebq�W3.1���_	�W�Ш��2I��v�k#�7@^�%�,�m5�:��ު�@9�ya&0h�\T�r��t.e㳚�Ql]!@�oJt�P��'�
7>NU��W飯�۫삘pvζ�������-}�.��.9'1���')�H����-ޕ�*<\&���<J��3�3��Xl��O���XB�5JJ�#]��Z�D�m��0q�\��P�yY�L/`s�E��kz�٨�$�i�~yҌuٸn�\�Q�l�ct��]��ֿ˘`��] X��a
�����b.x5� b/��չ�^8B�%w_�S�Jc��iL�3�K<�b���l6��+c�ڎu�KHf,�����"��;����mT˭$��HN���B"�o��}��A.팗b۫,��򒹤����}Dʤn �_yS;څ4��Y�(�OU�Ն�����w��k���W�E��5s�h#E�����D~L���U�ۦ�Q���.@�u;���_��o^D��G�Ov�;.F��jG�c�y!+��GO��!�vĆY�f��Ꮜ�df�4��vL�DI���b�����M�!Cm�ȅ!��t=U���6��Ox�ɼ{9�F��GV_<)w���7B6o�٩׷�f|VC0e�|Q�[���t�D�c�M�z�AC[q��i���p�u�{���r6�i,��n��C2��Mm��n��x����][��al)kG�-��0m["��OZ�����"�O:��.۷0� �����[�7+��>�Ml@�c3t:��I�Dy��>��ex�=�@{87X��Zx~�#�K�B� �vV�nGn�4<Ԣ�2��� sW�pC��c����n�v���7Ͼ�3SvXwZ�~æ�gM�!����c�6`�6����:*x%���sw:t��������#<ն��l������uLdW^��?��7�s��y���W����ǵ���8���l����\:�;��V�߂��)�̓���&���9r���6��b(�ޤ�H�'\���ؒ�����q�y�:�>;ؠ��X��ӅP��l�^����nun=:�����?-���]���7�~U�яC��ë�e|e��u�{��=ƞ#��]����f�/�wt��-������U�?�r�<%�GP4ٻoB߮n�p�Vvs�nأQa�bҏu�#BC����f���z�'Р�%��#����<���1�֕�PG���}�W��I��(��ƅ���M��M`��� �;��J�,��k�ߘN{,e@T�g
�/��n���p8�*�V��hI��}(��B�H�l܅qن��:)͋��d>x1��+m��>�RBa.�q@	�3߹���w�̜d>������Lo�1�Y�HVސ�y�D�D�Gnj��T?ҾAh�4+�2�[�s�ʖ�oq��b`br��O.s!�\�o��j���Sb�-�YE�M����a�κ˻�����\����4cV���4�-K|�ܴ;�81�d7����p�e�a�^��r:�u_��{WU��DamM"-6�y���@�@���`� eO3�����p����.�,�.��-[ذ�g��DpJ�$��!��k1��q�.<.��Y����k��u���QwJ�K��.���©���W8������$9GxNJ Z��4;���t4�K6v����\��Z���d�Tr�̯��bH�������}�b�����㧸���u�R47f\��Q��en�@��D��<��N�47��IP*���^��М~�-� ��7���)�C�ԧA2&~�eV�����WM�#0i�È=5J;	��t��1d�$�"T
���)�2p���".+�Ľ2(���o�
e���C�I}��|�Ob��$\`x CA�0AK��WS��k^CfWn��k�X�8��ç�.���ZP���~{�x�������q��xBH�����;����i�7PX_�Ī�bZ%mӠ_ŗ�!3ү
�`]�E��P�����:a�X�� �VMإ���3gvbamer4B|qo�N���)�iE�M���fKjz�-̑920k�&<��Z�R��Eq�l<u��Ju��F���<����j`�q��z�#�,�?�t<�LA��!Y�ǯ��K~ttOB�ʱ/�Zo�����癝C.����J)E?�p
�u^����-���Ŝ>�䟎g�"�1L�w��7����G���*��+:��!�Yu^���h\! F��0��{�%�X�o`��~8V|Z.׬:f��#��{�.
[��"��oc*��eL��D�%^�G���t�����?�d��$1�|��!p퍄ճn��@��H�t�q�&mǰ��$��[$8ǈA4�)	�t*3���=�)yp��En?�E�8��Q[�<:�-�:*�PSud��I ��-��V*-E��U�uq�k6\P��6L������Ҹ��\��n�!Zr�^�А@0�	��;E��-�{�x�M~�{/ԙk�6�[3��u���� ���9~��]��z��Xia�9G�E�l�w�!m�vV:ce�p�\�2�{,�'�X&�[����݁��Ƽ���SQ�|�{�� ������(}���8�����ڀ[�J����8^+�+���_�i!�������}_X���^P)��e��1[8�͂���^�������GLd�^#�H����I��%|-	��aֺ�$Z��n_��G��� !q�F���>N�:t�L������K��܀R���Q+yS��G+3pc�Z�\�W�	��ZСf��(���Jq��0H�p�Ԝ�o*掭B�ޣ*�kc���#��Q&.���E�zu-ތ�Z��=!�e�]�l_�{�E�T*J<n�Wn4�A(S&���~������8�i��"��Γ��5��֪0$)���G&o6�.��$�!��������!��d���/s�`��'�C-�Xy6���f��zҬ�����[�)�\\G̀�՗�}d�g��Tn�������]t��Q7ԕ�� Du��F��_��ь�2,;�ȋ�o���oC��)V�}�>q�{�Wx)|)Y���{>�N��s�����/=�7C13�^q�N����ϔ�(��a�=gsx�2��:S���va���t�d�:c��8��z#�w�R�_�� 45�$%R@����#A���vE\ʖ�����m˖H�{(f�h-�"��h=�`�"ؚ����XQ}�U�.�#)}R��t���&q�� �/����PZ�5N��w���1]��9���C���S��C+m0�Jz%�Xx�}I?�-ϙvR_J~^+�I�fI� �L�y���k�=�`