XlxV61EB    1f39     790 ��do�Ż�t�-|�r|��B��) �59{nJ�>E��4�w���%)A
6�T���/C�#S�~ߕ��ѭ�)�3c�n��$�;��ĥʧ	�]�u%g�B(Ԛ�"ㅊ&��ܐ%65�qX�g�b��Z��\L���;��,R���}L�i����ұk�L˕����~����<��X�7F����<�k=��w� ���-���J���!��kT�6â��Zv�z?��xu���k̔uÊi��Y�(�2ќ��5�?�'=dz6Ğ��'j{k�V-���(�a�"�A����Oo&嫜�$�9/����Z]��H��}������Y���g��d�kň� �TǠH�c�^�0���D�h�Д��'7 ��[E�}=��.��AJmӼo�r�]Og��-d %�އ�d���j1I����������H���r&A��7�M*or�GP����P�fݺ+�ʽ�Iя8&�`d9{KŃ��4��0���8�l��{�G~�m��ib����#�+j	)Z�a=�#��RC�
y.sY����wQ�3�b΢+�&��6_ lE�~�����Pd�QJ�f"o���`0�B�̂変��bsH�$en,�A�,�31�2�Y���f�G/�ؖ�)�z�� ��RskѣtS��>)�|�Ke�4�MȷG�aӭ�����?r��hNa�{)��wn�z0�8Y٫'(9:ӂ���MɚZ܃6��y����8�?�c�w���h=��ј�ǼT`\ʇc?��z�C'\�<T�ڞ�_��L�d>0ϗs�k4p�:՝A�l��k4��vM�	Ny_uk�;�c碊'��0�)<��r��3��ٍ��MD��G��{~BI���r���_�B���q��u�VC<�^~TZ3�b��73�hfA�k'z�g�����"b�0�t;=Rk� �#�3}�x
����W
�Y�>5�B��eX:C ���A�y�p�g[1��ӹ�C���	cP��dvs%�u&L������	�(�E�P��[c��G�mIsؿ���\g��2�l�k��󐧡����eAyls����*�C�Ӧ�N��0.�^�f�g��QWNBy�8/��z?TV��7��06��y$�n=�e\�<�U���b����Ni���+����^�Pn�B���zU��´�3g�l%��%#$�9��
.�?�OF��"�q�?*�I����Z`�u0p���o*��s��.��D���{{����5:&���d���zQO�Ȩ֕�=.e�ne<�A�Do��X����1��.�^�y����tQ���)��K1��V3u. �0K�u0�:q�
B���3�+�ߩ.��{x�M���)^.w�G����0��5�)0muKr�y�!�_�-P(B��T�^9��D��7���ݤ�4����S.5nW�&Ln/2���z6w��@e�!(��},��P���OF�EO���!��M�����%������:2����0��3�ܯCu��c����u �+�ѷ�g���%8@t���:}���@�;������؇�3�*ƅy"fz���X������/^��_���tK��a��7���.�`��~�\R2�y�=r�USђ~]�~=�'�M�=�� �w J��	K�<^
��=X0���?�6'�f/z�9��ӎ��Bn��|3�+ò���x�������5��墒�q?��oyё��a�U��fP}���ٕ��黫�)	t�&�p�����������P�_\�V 'ȗ]�JZ@�B��-��e
Vd1�u��:R*91޺p���2���;>m����[�O���vK�/b����� �قE�ݑzx�$�B��%����j�өX)�'v��#����K��Y�up�� y2cet�-V+`��d0��rB�Y��LY�a|�