XlxV61EB     647     180r+�9 �#�Q�"$���'깹u�K�[�ܜcX�=U7������ݍT#�S��X��lMF�׈ŤȻLE&5c�O\y���5nOa�hf���mv�Na�- ��	�&��BO�%:�P�/���Uj�t:P
�x�^���Tr7��|�o���{����}v2%M�eO��-E�������k�A�I%��tT��h��<.�2���=:0��}��5�9*�������S�����&�
s��m�]5/l�}ԨS��U�4�i�t���H��g�s���]����O2bQ�U�7��^�+���G>B2.��^�:
p'�l��ٓ�p�)@�����Cx��wQJNM�S�Ai�ӫ=�V+2�F	���l�]